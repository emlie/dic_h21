// Module for the 2 x 2 pixel array using pixelSensor

// Include the pixel sensor files
`include "pixelSensor.fl";

// Use the pixel sensor in the pixel array
//
// Signals that need to be in a bus:
// - DATA
//
// Signals that are common for the pixels
// -
module pixelArray (
    ports
);
    
endmodule